interface sr_interface(input clk, rst);
  logic [4:0] addr;
  logic [15:0] din;
  logic wr_en;
  logic [15:0] dout;
  
  
  
endinterface
  
  